`timescale 1ns/1ps
module simple(
    input wire clk_i
);
endmodule
