`ifndef ALU_PKG_SV
`define ALU_PKG_SV

`timescale 1ps/1ps
package alu_pkg;
  typedef enum logic[3:0] {
    ALU_ADD  = 4'b0000,
    ALU_SUB  = 4'b0001,
    ALU_AND  = 4'b0010,
    ALU_OR   = 4'b0011,
    ALU_XOR  = 4'b0100,
    ALU_SLT  = 4'b0101,
    ALU_SLTU = 4'b0110,
    ALU_SLL  = 4'b0111,
    ALU_SRL  = 4'b1000,
    ALU_SRA  = 4'b1001
  } alu_op_e;

  typedef enum logic[1:0] {
    ALU_SRC_REG     = 2'b00,  // Register
    ALU_SRC_IMM     = 2'b01,  // Immediate
    ALU_SRC_PC      = 2'b10,  // PC (for AUIPC)
    ALU_SRC_FOUR    = 2'b11   // Constant 4 (for JAL/JALR)
  } alu_src_e;

endpackage

`endif // ALU_PKG_SV
